��  CCircuit��  CSerializeHack           ��  CPart              ���  CLED_Y�� 	 CTerminal  ���     
   ����`�?	5\��?;  
�  ���        "��`�?	5\��?�    ����         ����    ��  CChain��  CRotateKnob  ����          5    7 �  ����         � V  y 7 �� 	 CMechTerm@�z�P�@      ��        y 7 �   �@�z�P�@      ��        y 7 @ p   � ]    ����     	 @�z�P�@                    pu     	 @�z�P�@          �0\t<�@      Ľ         7 P   �0\t<�@      ĽUUUUUUN� 7   P    $    `�e�     	 0\t<�@UUUUUUN�            �p�u     	 0\t<�@              dt�         P�    p   8J��=>0\t<�@Y
!Q6��?� `f����1;Zx>@�z�P�@�6$��? 3���<  ��7 p       5         y @ 7 p      � V &       0\t<�@Y
!Q6��?@�z�P�@�6$��?��  CMotorEM
�  �	�           ~�`�?����>4�<  
�  	        "��`�?����>4��  �0\t<�@      Ľ    �P�                  ��     	 0\t<�@    �P�    ��        ��      bK�6�>0\t<�@�*�����?��̘�gr�0\t<�@�*�����?��  CSPST��  CToggle  �� ��         
�  ��1       ?D0K
 "@          
�  ��1     	   I���`�?            �� �          ����P    �� 	 CResistor��  CDummyValue  8(8(    680           @�@      �?   
�  ((=)     	   I���`�?          
�  t(�)        I���`�?            <!t1     &      ��8 	  ��  CLED
�  ��1        I���`�?����N�;  
�  ��1          ~�`�?����N��    �� �     *    ����    ��  �P�t      ,  
�  ����       ?D0K
 "@          
�  ����     
   ����`�?            �r��     .    ����P    "�$�  @�@�    680           @�@      �?   
�  0�E�     
   ����`�?�����ۛ�  
�  |���        ���`�?�����ۛ;    D�|�     2      ��8 	  ��  CLED_G
�  ����        ���`�?ߔ=i���  
�  ����          ~�`�?ߔ=i��;    �d��     6    ����    �� 
 CBattery9V$�  �p�p    9V            "@      �? V 
�  �`�u           ~�`�?x�in��  
�  �`�u        ?D0K
 "@�M4�s�)=    tt�      ;    ��   �  ��  CBuzzer
�  �� ��       	   I���`�?�D����<  
�  �L�a          ~�`�?�D�����    T� �L     ?    ��  6 `  "�$�  @@    680           @�@      �?   
�  0E     
   ����`�?oooo���<  
�  |�        "��`�?oooo����    D|!     C      ��8 	                ���  CWire  �	      F�  ��      F�  � �       F�   1     
 F�  �!     
 F�    !      
 F�    �     
 F�  ����      F�  �(�)      F�  � ��      	 F�  @�a�     F��� 
 CCrossOver  .�4�    ��  �A�     F�  �1�      F�  ��	�      F�  �	�       F�  0)1     	 F�  � 	1      	 F�  0�1�      
 F�  (()1      	 F�  �(�1       F�  �0�1      F�   0�1      F�   `�a      F�   �!a       F�   ���      F�   0!�       F�   p1q      F�   `q       F�  �`a      F�  �0	1     	 F�  0`�a      F�  �011      F�  001a       F�  0`1�       F�S�  .�4�    ��  0�1q       F�  ���      
 F�  ����     
 F�  ��1�     
               �                              M   I          Q       W    G   R     ^ ! ! f & [ & ' ' O * * ] + + h . . a / / n 2 Z 2 3 3 N 6 6 N 7 7 V ; e ; < _ < ? P ? @ @ g C J C D D H H  D I  G K C m L M J L  3 6 ' \ Y ? R  R l  Q V k 7 W U  f [ P X 2 o & X O ] \ * b   ` < b _ ` . ^ a d k e c ; d ! Y j @ + i h g i U k T j c o K / m n Z            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 